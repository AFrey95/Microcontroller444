library verilog;
use verilog.vl_types.all;
entity test_file is
end test_file;

library verilog;
use verilog.vl_types.all;
entity test_controller is
end test_controller;

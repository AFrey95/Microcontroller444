library verilog;
use verilog.vl_types.all;
entity altsyncram is
    generic(
        address_aclr_a  : string  := "UNUSED";
        address_aclr_b  : string  := "NONE";
        address_reg_b   : string  := "CLOCK1";
        byte_size       : integer := 8;
        byteena_aclr_a  : string  := "UNUSED";
        byteena_aclr_b  : string  := "NONE";
        byteena_reg_b   : string  := "CLOCK1";
        clock_enable_input_a: string  := "NORMAL";
        clock_enable_input_b: string  := "NORMAL";
        clock_enable_output_a: string  := "NORMAL";
        clock_enable_output_b: string  := "NORMAL";
        indata_aclr_a   : string  := "UNUSED";
        indata_aclr_b   : string  := "NONE";
        indata_reg_b    : string  := "CLOCK1";
        init_file       : string  := "UNUSED";
        init_file_layout: string  := "PORT_A";
        intended_device_family: string  := "UNUSED";
        implement_in_les: string  := "OFF";
        lpm_hint        : string  := "UNUSED";
        lpm_type        : string  := "altsyncram";
        maximum_depth   : integer := 0;
        numwords_a      : integer := 0;
        numwords_b      : integer := 0;
        operation_mode  : string  := "BIDIR_DUAL_PORT";
        outdata_aclr_a  : string  := "NONE";
        outdata_aclr_b  : string  := "NONE";
        outdata_reg_a   : string  := "UNREGISTERED";
        outdata_reg_b   : string  := "UNREGISTERED";
        power_up_uninitialized: string  := "FALSE";
        ram_block_type  : string  := "AUTO";
        rdcontrol_aclr_b: string  := "NONE";
        rdcontrol_reg_b : string  := "CLOCK1";
        read_during_write_mode_mixed_ports: string  := "DONT_CARE";
        width_a         : integer := 1;
        width_b         : integer := 1;
        width_byteena_a : integer := 1;
        width_byteena_b : integer := 1;
        widthad_a       : integer := 1;
        widthad_b       : integer := 1;
        wrcontrol_aclr_a: string  := "UNUSED";
        wrcontrol_aclr_b: string  := "NONE";
        wrcontrol_wraddress_reg_b: string  := "CLOCK1";
        clock_enable_core_a: string  := "USE_INPUT_CLKEN";
        clock_enable_core_b: string  := "USE_INPUT_CLKEN";
        enable_ecc      : string  := "FALSE";
        read_during_write_mode_port_a: string  := "NEW_DATA_NO_NBE_READ";
        read_during_write_mode_port_b: string  := "NEW_DATA_NO_NBE_READ"
    );
    port(
        wren_a          : in     vl_logic;
        wren_b          : in     vl_logic;
        rden_a          : in     vl_logic;
        rden_b          : in     vl_logic;
        data_a          : in     vl_logic_vector;
        data_b          : in     vl_logic_vector;
        address_a       : in     vl_logic_vector;
        address_b       : in     vl_logic_vector;
        clock0          : in     vl_logic;
        clock1          : in     vl_logic;
        clocken0        : in     vl_logic;
        clocken1        : in     vl_logic;
        clocken2        : in     vl_logic;
        clocken3        : in     vl_logic;
        aclr0           : in     vl_logic;
        aclr1           : in     vl_logic;
        byteena_a       : in     vl_logic_vector;
        byteena_b       : in     vl_logic_vector;
        addressstall_a  : in     vl_logic;
        addressstall_b  : in     vl_logic;
        eccstatus       : out    vl_logic_vector(2 downto 0);
        q_a             : out    vl_logic_vector;
        q_b             : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of address_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of address_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of address_reg_b : constant is 1;
    attribute mti_svvh_generic_type of byte_size : constant is 1;
    attribute mti_svvh_generic_type of byteena_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of byteena_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of byteena_reg_b : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_input_a : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_input_b : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_output_a : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_output_b : constant is 1;
    attribute mti_svvh_generic_type of indata_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of indata_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of indata_reg_b : constant is 1;
    attribute mti_svvh_generic_type of init_file : constant is 1;
    attribute mti_svvh_generic_type of init_file_layout : constant is 1;
    attribute mti_svvh_generic_type of intended_device_family : constant is 1;
    attribute mti_svvh_generic_type of implement_in_les : constant is 1;
    attribute mti_svvh_generic_type of lpm_hint : constant is 1;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of maximum_depth : constant is 1;
    attribute mti_svvh_generic_type of numwords_a : constant is 1;
    attribute mti_svvh_generic_type of numwords_b : constant is 1;
    attribute mti_svvh_generic_type of operation_mode : constant is 1;
    attribute mti_svvh_generic_type of outdata_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of outdata_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of outdata_reg_a : constant is 1;
    attribute mti_svvh_generic_type of outdata_reg_b : constant is 1;
    attribute mti_svvh_generic_type of power_up_uninitialized : constant is 1;
    attribute mti_svvh_generic_type of ram_block_type : constant is 1;
    attribute mti_svvh_generic_type of rdcontrol_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of rdcontrol_reg_b : constant is 1;
    attribute mti_svvh_generic_type of read_during_write_mode_mixed_ports : constant is 1;
    attribute mti_svvh_generic_type of width_a : constant is 1;
    attribute mti_svvh_generic_type of width_b : constant is 1;
    attribute mti_svvh_generic_type of width_byteena_a : constant is 1;
    attribute mti_svvh_generic_type of width_byteena_b : constant is 1;
    attribute mti_svvh_generic_type of widthad_a : constant is 1;
    attribute mti_svvh_generic_type of widthad_b : constant is 1;
    attribute mti_svvh_generic_type of wrcontrol_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of wrcontrol_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of wrcontrol_wraddress_reg_b : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_core_a : constant is 1;
    attribute mti_svvh_generic_type of clock_enable_core_b : constant is 1;
    attribute mti_svvh_generic_type of enable_ecc : constant is 1;
    attribute mti_svvh_generic_type of read_during_write_mode_port_a : constant is 1;
    attribute mti_svvh_generic_type of read_during_write_mode_port_b : constant is 1;
end altsyncram;
